`timescale 1ns/1ps

module I2C_TB;
    reg [6:0] Address;
    reg [7:0] Data_Frames;
    reg rw;
    reg processor;
    reg writes;

    wire [3:0] shtreads, bytesreceived, outputreceivedcounter;
    wire [2:0] masterstateout;
    wire [7:0] datareceived;
    wire [15:0] tempoutput, rhoutput;
    wire [2:0] sclstateout;
    
    clock_gen testclk1 (clk);

    shtack testack (
        .clk (clk),
        .Master_State_Out(masterstateout),
        .Sda_Data(Sda_Data),
        .Scl_Data(Scl_Data)
        );
    
    i2c_master master1 (
        .clk (clk), 
        .Sda_Data(Sda_Data), 
        .Processor_Ready(processor), 
        .Command_Data_Frames(Data_Frames),
        .Peripheral_Address(Address),
        .Scl_Data(Scl_Data),
        .i2c_writes(writes),
        .SHT_Reads(shtreads),
        .CRC_Error(CRC_Error),
        .Bytes_Received(bytesreceived),
        .Data_Received(datareceived),
        .Output_Received_Counter(outputreceivedcounter),
        .Frames_Read(Frames_Read),
        .Master_State_Out(masterstateout),
        .r_or_w(rw),
        .Scl_State_Out(sclstateout)
        
        );
    i2c_sht40 peripheral1 (
        .clk (clk),
        .Output_Received_Counter(outputreceivedcounter), 
        .Data_Received(datareceived), 
        .SHT_Reads(shtreads), 
        .Temperature_Output(tempoutput), 
        .Humidity_Output(rhoutput),
        .Temp_Ready_Out(Temp_Ready_Out),
        .RH_Ready_Out(RH_Ready_Out)
        );
    i2c_scl scl1 (
        .clk(clk),
        .Scl_Data(Scl_Data),
        .Sda_Data(Sda_Data),
        .Master_State_Out(masterstateout),
        .Scl_State_Out(sclstateout)
    );

    initial begin
        Address = 7'b1000100; //0x44 in hex
        Data_Frames = 8'b11111101; //0xfd in hex
        rw = 1'b0;
        processor = 1'b1;
        writes = 1'b1;
    end
    
    pullup SCL (Scl_Data);
    pullup SDA (Sda_Data);

endmodule

module clock_gen (output reg clk);
    initial begin
        clk = 0;
    end
    
    always begin
        #1 clk = ~clk;
        
    end
endmodule

module shtack (input clk, inout Sda_Data, input [2:0] Master_State_Out, input Scl_Data);
    reg sdadatalocal;
    reg sdaflag; 
    reg scledgechecker;
    reg [3:0] Counter; 

    initial begin
        sdadatalocal = 1'bZ;
        scledgechecker = 1'b0;
        Counter = 4'd0;
    end

    assign Sda_Data = sdadatalocal;

    always @(posedge clk) begin
        if (Master_State_Out == 3'b010 || Master_State_Out == 3'b100 || Counter > 4'd7) begin
            scledgechecker <= Scl_Data;
            if (scledgechecker && ~Scl_Data) begin
                Counter <= Counter + 4'd1;
            end 
            if (Counter == 4'd8) begin
                sdadatalocal <= 1'b0; 
            end
            if (Counter == 4'd9) begin
                sdadatalocal <= 1'bZ;
                Counter <= 4'd0;
            end
                   
        end
    end 
endmodule